module arbiter(
    input logic clk,
    input logic rst,
    input logic [255:0] arb_mem_req,
    output logic [255:0] arb_mem_resp
);



endmodule : arbiter