import rv32i_types::*;

module MEM_WB(


);




endmodule : MEM_WB