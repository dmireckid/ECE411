import rv32i_types::*;

module ID(


);



endmodule : ID