import rv32i_types::*;

module cpu(



);


endmodule : cpu