import rv32i_types::*;

module ID_EX(
    input clk,
    input rst,
    input pc_out_IFID,
    output rv32i_word pc_out_IDEX,
    //figure out instruction stuff

);




endmodule : ID_EX