import rv32i_types::*;

module WB(


);




endmodule : WB