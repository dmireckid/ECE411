import rv32i_types::*;

module IF(


);


endmodule : IF