import rv32i_types::*;

module mp3(





);










endmodule : mp3