import rv32i_types::*;

module IF_ID(


);




endmodule : IF_ID