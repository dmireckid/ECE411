import rv32i_types::*;

module MEM(


);



endmodule : MEM