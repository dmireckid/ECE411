import rv32i_types::*;

module ID_EX(


);




endmodule : ID_EX