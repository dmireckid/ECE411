import rv32i_types::*;

module control_rom(



);




endmodule : control_rom