import rv32i_types::*;

module MEM(
    input clk,
    input rst,
    input rv32i_word inst,
    input rv32i_word pc_in,
    input rv32i_word rs1_in,
    input rv32i_word rs2_in,
    input rv32i_control_world MEM_ctrl_in,



);

    



endmodule : MEM